module uart_rx (
    input clk,
    input reset,
    input rx_data,
    output reg [15:0] data_out
);

// Implement UART receiver logic to buffer received data
// and output a 16-bit value when a complete word is received

endmodule
